//-----------------------------------------------------------------------
// Author : Golovachenko Victor
//-----------------------------------------------------------------------
`define C_I2C_MASTER_CORE_IDLE     3'h0
`define C_I2C_MASTER_CORE_START    3'h1
`define C_I2C_MASTER_CORE_RESTART  3'h2
`define C_I2C_MASTER_CORE_STOP     3'h3
`define C_I2C_MASTER_CORE_TXBYTE   3'h4
`define C_I2C_MASTER_CORE_RXBYTE   3'h5
